//
/* 
    multi-line comment.  Uses a nested lexer.  Is there a way to drop back
    rather than recurse into?
*/
 
module hello1(a,b,f,d);

endmodule

module hello2(a,b,f,d);

    parameter p = 1'b1 + 10'd2 / 4;
    parameter d = f;
    
    input a;

endmodule



